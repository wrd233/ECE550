module not_gate(
  input a,
  output out
);
  not my_and(out,a);
endmodule
