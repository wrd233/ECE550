module alu(data_operandA, data_operandB, ctrl_ALUopcode, ctrl_shiftamt, data_result, isNotEqual, isLessThan, overflow);

    input [31:0] data_operandA, data_operandB;
    input [4:0] ctrl_ALUopcode, ctrl_shiftamt;

    output [31:0] data_result;
    output isNotEqual, isLessThan, overflow;

//    // YOUR CODE HERE //
//    always @(ctrl_ALUopcode, data_operandA, data_operandB) begin
//        case(ctrl_ALUopcode)
//            // TODO: 根据情况调用函数
//            0:  // ADD
//            1:  // SUBTRACT
//            2:  // AND
//            3:  // OR
//            4:  // SLL
//            5:  // SRA
//        endcase
//    end
endmodule
