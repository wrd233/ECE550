module or_gate(
  input a,
  input b,
  output out
);
  or my_and(out,a,b);
endmodule
