module and_gate(
  input a,
  input b,
  output out
);
  and my_and(out,a,b);
endmodule
