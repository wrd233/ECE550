module nor_gate(
  input a,
  input b,
  output out
);
  nor my_norg(out,a,b);
endmodule
