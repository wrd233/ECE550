module alu_1_bit;

endmodule
